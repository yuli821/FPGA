//-------------------------------------------------------------------------
//      ECE 385 - Summer 2021 Lab 7 Top-level                            --
//                                                                       --
//      Updated Fall 2021 as Lab 7                                       --
//      For use with ECE 385                                             --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module game (

      ///////// Clocks /////////
      input    MAX10_CLK1_50,

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,





      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);

//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
	logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0, score; //4 bit input hex digits
	logic [1:0] signs;
	logic [1:0] hundreds;
	logic [7:0] keycode [6];
	logic key[10];
	logic i2c_serial_scl_in, i2c_serial_scl_oe, i2c_serial_sda_in, i2c_serial_sda_oe;
	logic [1:0] aud_mclk_ctr;
	logic [15:0] audio_data;
	logic [13:0] audio_address;
	logic count_en;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ;
	assign USB_IRQ = ARDUINO_IO[9];
	
	//Assignments specific to Sparkfun USBHostShield-v13
	//assign ARDUINO_IO[7] = USB_RST;
	//assign ARDUINO_IO[8] = 1'bZ;
	//assign USB_GPX = ARDUINO_IO[8];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[8] = 1'bZ;
	//GPX is unconnected to shield, not needed for standard USB host - set to 0 to prevent interrupt
	assign USB_GPX = 1'b0;
	
	//HEX drivers to convert numbers to HEX output
	HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
	assign HEX4[7] = 1'b1;
	
	HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
	assign HEX3[7] = 1'b1;
	
	HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
	assign HEX1[7] = 1'b1;
	
	HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
	assign HEX0[7] = 1'b1;
	
	//fill in the hundreds digit as well as the negative sign
	//assign HEX5 = {1'b1, ~signs[1], 3'b111, ~hundreds[1], ~hundreds[1], 1'b1};
	HexDriver hex_driver5 (score, HEX5[6:0]);
	assign HEX5[7] = 1'b1;
	
	assign HEX2 = {1'b1, ~signs[0], 3'b111, ~hundreds[0], ~hundreds[0], 1'b1};
	
	
	assign {Reset_h}=~ (KEY[0]); 
	
	assign i2c_serial_scl_in = ARDUINO_IO[15];
	assign ARDUINO_IO[15] = i2c_serial_scl_oe ? 1'b0 : 1'bz;
		
	assign i2c_serial_sda_in = ARDUINO_IO[14];
	assign ARDUINO_IO[14] = i2c_serial_sda_oe ? 1'b0 : 1'bz;
	
	assign ARDUINO_IO[1] = ARDUINO_IO[2];
//	assign ARDUINO_IO[2] = ARDUINO_IO[1];
//	assign ARDUINO_IO[1] = 1'bz;

	assign count_en = (key[2]||key[6]);  //test
	
	assign ARDUINO_IO[3] = aud_mclk_ctr[1];
	//generate 12.5 MHz CODEC mclk
	always_ff @ (posedge MAX10_CLK1_50) begin
			aud_mclk_ctr <= aud_mclk_ctr + 1'b1;
	end

	
	//remember to rename the SOC as necessary
	game_soc u0 (
		.clk_clk                           (MAX10_CLK1_50),    //clk.clk
		.reset_reset_n                     (1'b1),             //reset.reset_n
		.altpll_0_locked_conduit_export    (),    			   //altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (), 				   //altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),     			   //altpll_0_areset_conduit.export
    
		.key_external_connection_export    (KEY),    		   //key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),            				   //clk_sdram.clk
	   .sdram_wire_addr(DRAM_ADDR),               			   //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                			   //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),              		   //.cas_n
		.sdram_wire_cke(DRAM_CKE),                 			   //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                		   //.cs_n
		.sdram_wire_dq(DRAM_DQ),                  			   //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),                //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),              		   //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                		   //.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.hex_digits_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),
		.leds_export({hundreds, signs, LEDR}),
		.keycode0_export({keycode[2],keycode[1],keycode[0]}),
		.keycode1_export({keycode[5],keycode[4],keycode[3]}),
		
		.i2c0_sda_in(i2c_serial_sda_in),
		.i2c0_scl_in(i2c_serial_scl_in),
		.i2c0_sda_oe(i2c_serial_sda_oe),
		.i2c0_scl_oe(i2c_serial_scl_oe)
//		
	 );
	 //A:0 D:1 W:2 F:3 <-:4 ->:5 up:6 sp:7 en:8 esc:9
	 vga_sprite_controller v0(.CLK(MAX10_CLK1_50), .RESET(Reset_h), .key(key),
					.red(VGA_R), .green(VGA_G), .blue(VGA_B), .hs(VGA_HS), .vs(VGA_VS),
					.score(score));
					
	 keycode_reader key0(.keycode(keycode), .key(key));
	 
	 counter c0(.Reset(Reset_h), .Clk(ARDUINO_IO[4]), .en(count_en), .address(audio_address));
		
	 //audio_ram ram0(.address(audio_address), .clock(ARDUINO_IO[4]), .q(audio_data));
	 RAM_audio (.data_In(), .write_address(),.read_address(audio_address),.we(1'b0),
					.Clk(ARDUINO_IO[5]),.data_Out(audio_data));
		
	 codec codec0(.sample({audio_data,8'b0}), .SCLK(ARDUINO_IO[5]), 
						.LRCLK(ARDUINO_IO[4]), .Reset(Reset_h), .out(ARDUINO_IO[2]));
	 

endmodule
