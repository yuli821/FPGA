module tile_rom(output logic [0:29][0:39] Tile);
						
		
		assign Tile = ROM;
		
		parameter [0:29][0:39] ROM = 
		{
		40'hFFFFFFFFFF, // will occupy about two line if not zero. HOW COME?!!!!
		40'h8000000001, // 1
		40'h8000000001, // 2
		40'h8000000001, // 3
		40'h81FF000001, // 4
		40'hC003000001, // 5
		40'h8000FFFFFF, // 6
		40'h8000000001, // 7
		40'hFF00000001, // 8
		40'h8080000001, // 9
		40'h8000000001, // 10
		40'h8000000001, // 11
		40'hFFFFFFFFE1, // 12
		40'h80000003E1, // 13
		40'h8000000001, // 14
		40'h8000000001, // 15
		40'h8CFFFFF001, // 16
		40'h8000003FFF, // 17
		40'h8000000001, // 18
		40'h8000000001, // 19
		40'h8000000001, // 20
		40'hFFFFFE0001, // 21
		40'h8000008001, // 22
		40'h800000FFC1, // 23
		40'h8000000001, // 24
		40'hFFFFF00001, // 25
		40'h800000000F, // 26
		40'h8000000001, // 27
		40'h8000000001, // 28
		40'hFFFFFFFFFF  // 29
		};

		
endmodule

		